

module test;
  int mat[3][3] = '{ '{1,2,3},'{4,5,6},'{7,8,9} };
  int t;

  initial begin
    $display("%p",mat);
        
     
  end


endmodule


//  1 2 3
//  4 5 6
//  7 8 9
//
//  7 8 9 
//  4 5 6 
//  1 2 3
//
//  7 4 1
//  8 5 2
//  9 6 3
