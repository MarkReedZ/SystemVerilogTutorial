

module block( input clk, reset_n,push,pop,valid,ready,ack,x,y,xone,xtwo );
  logic test;
endmodule


