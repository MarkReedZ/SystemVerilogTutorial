
timeskew checks peterfab.com specify block
