
interface valid_intf (/*AUTOARG*/
   );
input logic             clk;
input logic             reset_n;
input logic             valid;
input logic             ack;

endinterface

