
module hello;
  int x;

  initial begin

    $display("Hello World. x is %0d", x);

  end

endmodule

