
module test;
  /* my_intf AUTO_TEMPLATE "\(.*\)_my_i" (
      .clk       (clk_@),
      .reset_n   (reset_n_@),
      .\(.*\)    (),
  )*/
  
  my_intf a_my_i ( /*AUTOINST*/ );
  my_intf b_my_i ( /*AUTOINST*/ );

endmodule
